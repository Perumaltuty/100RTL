`timescale 1ns / 1ps
module buffer(a,y);
	input a;
	output y;
	assign y=a;	
endmodule
