module clock_freq(clock);
input clock;
endmodule
